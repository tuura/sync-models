module Untitled (n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29);
    
    output n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
    
    INV b0 (.I(n0), .ON(n1));
    BUF b1 (.I(n1), .O(n2));
    BUF b2 (.I(n2), .O(n3));
    BUF b3 (.I(n3), .O(n4));
    BUF b4 (.I(n4), .O(n5));
    BUF b5 (.I(n5), .O(n6));
    BUF b6 (.I(n6), .O(n7));
    BUF b7 (.I(n7), .O(n8));
    BUF b8 (.I(n8), .O(n9));
    BUF b9 (.I(n9), .O(n10));
    BUF b10 (.I(n10), .O(n11));
    BUF b11 (.I(n11), .O(n12));
    BUF b12 (.I(n12), .O(n13));
    BUF b13 (.I(n13), .O(n14));
    BUF b14 (.I(n14), .O(n15));
    BUF b15 (.I(n15), .O(n16));
    BUF b16 (.I(n16), .O(n17));
    BUF b17 (.I(n17), .O(n18));
    BUF b18 (.I(n18), .O(n19));
    BUF b19 (.I(n19), .O(n20));
    BUF b20 (.I(n20), .O(n21));
    BUF b21 (.I(n21), .O(n22));
    BUF b22 (.I(n22), .O(n23));
    BUF b23 (.I(n23), .O(n24));
    BUF b24 (.I(n24), .O(n25));
    BUF b25 (.I(n25), .O(n26));
    BUF b26 (.I(n26), .O(n27));
    BUF b27 (.I(n27), .O(n28));
    BUF b28 (.I(n28), .O(n29));
    BUF b29 (.I(n29), .O(n0));
    
    // signal values at the initial state:
    // !n0 !n1 !n2 !n3 !n4 !n5 !n6 !n7 !n8 !n9 !n10 !n11 !n12 !n13 !n14 !n15 !n16 !n17 !n18 !n19 !n20 !n21 !n22 !n23 !n24 !n25 !n26 !n27 !n28 !n29
    
endmodule
