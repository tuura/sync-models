module BUF_BUILTIN (output out, input inp);
    assign out = inp;
endmodule
