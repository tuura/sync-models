// vi: set ft=verilog :

{%- set ntransitions = nets|length %}

`define clk_rst @(posedge clk) disable iff (reset)

module spec (
          input reset
        , input clk
        , input [{{firebits-1}}:0] fire

        {%- for net in nets %}
        , input {{net}}
        {%- endfor %}

        {%- for net in nets %}
        , input {{net}}_precap
        {%- endfor %}

        {%- for output in stateless_outs %}
        , input {{ output }} // (stateless) output
        {%- endfor %}
    );

    {%- if ndbits %}

    reg {{ "[%d:0] " % (ndbits-1) if ndbits>1 -}} ndbits; // non-determinism bits
    {%- endif %}

    // fire signal constraints

    reg [{{firebits-1}}:0] fire_ne;  // fire, sampled on negedge

    always @(negedge clk)
        if (reset) fire_ne = 0; else fire_ne = fire;

    // Note:
    // - fire = [0, {{ntransitions-1}}] -> transition #fire is enabled
    // - fire = {{ntransitions}} -> no transitions enabled

    fire_in_range : assume property ( `clk_rst fire <= {{ntransitions}} );

    fire_cycle_stable : assume property(`clk_rst fire == fire_ne);

    // spec model

    integer state;

    always @(posedge clk or posedge reset) begin

        if (reset) begin

            {%- set initial_ind = state_inds[initial_spec] %}

            state <= {{ initial_ind }}; // {{ initial_spec }}

        end else begin
            {% for from, tr, to in transitions -%}
            {%- set signal     = tr[:-1]          -%}
            {%- set sign       = tr[-1]           -%}
            {%- set from_ind   = state_inds[from] -%}
            {%- set to_ind     = state_inds[to]   -%}
            {%- set verilog_tr = ("~" + signal) if sign == "-" else signal %}
            if (state == {{ from_ind }} && {{ verilog_tr }}) state <= {{ to_ind }};  // {{ to }}
            {%- endfor %}

        end

    end

    // Spec Compliance Properties:

    {%- for signal in inputs + outputs %}

    wire {{ signal }}_can_fall = 0
        {%- for prior, tr, _ in transitions if tr == signal + "-" %}
        {%- set prior_ind = state_inds[prior] %}
        {{ "|| (state == %d)"|format(prior_ind) }}
        {%- endfor -%}
        ;

    wire {{ signal }}_can_rise = 0
        {%- for prior, tr, _ in transitions if tr == signal + "+" %}
        {%- set prior_ind = state_inds[prior] %}
        {{ "|| (state == %d)"|format(prior_ind) }}
        {%- endfor -%}
        ;

    {%- endfor %}

    // Assumptions (spec compliance):
    {% for input in inputs %}
    compliance_{{input}}_rise: assume property ( `clk_rst $rose({{input}}) |-> {{input}}_can_rise );
    compliance_{{input}}_fall: assume property ( `clk_rst $fell({{input}}) |-> {{input}}_can_fall );
    {%- endfor %}

    // Assertions (spec compliance):
    {% for output in outputs %}
    compliance_{{output}}_rise: assert property ( `clk_rst $rose({{output}}) |-> {{output}}_can_rise );
    compliance_{{output}}_fall: assert property ( `clk_rst $fell({{output}}) |-> {{output}}_can_fall );
    {%- endfor %}

    // Enable signals:

    // Note: while internal transition enable status are indicated by (net ^
    // net_precap), inputs are generated by the environment and may therefore
    // may be enabled wile the expression (input ^ input_precap) is false.
    // Input enable status must therefore be derived from the spec, as
    // input_can_rise | input_can_fall.
    {% for input in inputs %}
    assign {{input}}_ena = {{input}}_can_rise | {{input}}_can_fall;
    {%- endfor -%}
    {%- for net in stateful_nets %}
    assign {{net}}_ena = {{net}}_precap ^ {{net}};
    {%- endfor %}

    // Output Persistency Properties:
    {% for net in stateful_nets %}
    persistency_{{net}}: assert property ( `clk_rst {{net}}_ena |=> ({{net}}_ena || ~$stable({{net}})) );
    {%- endfor %}

    // Deadlock

    // Deadlock freeness: on each cycle, at least one internal transition is
    // enabled or an input can change.

    assign exist_enabled_transition =
        {%- for input in inputs %}
        | {{input}}_ena
        {%- endfor -%}
        {%- for net in stateful_nets %}
        | {{net}}_ena
        {%- endfor -%}
    ;

    // For arbiter circuit:
    //
    // always_grant: assert property ( `clk_rst
    //     $rose(r1) |-> ##[1:$] ($rose(g1) | $rose(g2) | $rose(g3) | exist_enabled_transition)
    // );

    deadlock_free: assert property ( `clk_rst
        not (##[1:$] ~exist_enabled_transition)
    );

    // Transition firing assumptions: a transitions can only be fired when
    // it's enabled (i.e. when a stateful gate can capture a new value = its
    // input and output are different).

    {% for input in inputs %}
    {%- set pre_net = input + "_precap" %}
    {%- set fire_ind = loop.index0 -%}
    firing_{{fire_ind}}: assume property ( `clk_rst (fire == {{fire_ind}}) |-> ({{input}} ^ {{pre_net}}) );
    {% endfor -%}

    {% for net in stateful_nets %}
    {%- set fire_ind = loop.index0 + inputs|length -%}
    firing_{{fire_ind}}: assume property ( `clk_rst (fire == {{fire_ind}}) |-> ({{net}} ^ {{net}}_precap) );
    {% endfor %}
endmodule

module bind_info();

    bind circuit spec u1 (
          .reset(reset)
        , .clk(clk)
        , .fire(fire)

        {%- for net in nets %}
        , .{{net}}({{net}})
        {%- endfor -%}

        {%- for net in nets %}
        , .{{net}}_precap({{net}}_precap)
        {%- endfor -%}
    );

endmodule
