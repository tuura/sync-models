// vi: set ft=verilog :

{%- set inputs = spec["inputs"]|sort %}
{%- set outputs = spec["outputs"]|sort %}
{%- set initial = spec["initial_state"] %}
{%- set transitions = spec["transitions"]|sort %}
{%- set ntransitions = (inputs+stateful.values())|length %}

`define clk_rst @(posedge clk) disable iff (reset)

module spec (
          input reset
        , input clk
        , input [{{bit_size(ntransitions)-1}}:0] fire

        {%- for input in inputs %}
        , input {{ input }} // input
        , input {{ input }}_precap
        {%- endfor %}

        {%- for gate in stateful.values() %}
        , input {{ get_output_net(gate) }} // {{"output" if get_output_net(gate) in outputs else "internal"}}
        , input {{ get_output_net(gate) }}_precap
        {%- endfor %}

        {%- for output in stateless_outs %}
        , input {{ output }} // (stateless) output
        {%- endfor %}

    );

    {%- if ndbits %}

    reg {{ "[%d:0] " % (ndbits-1) if ndbits>1 -}} ndbits; // non-determinism bits
    {%- endif %}

    // fire signal constraints

    reg [{{bit_size(ntransitions)-1}}:0] fire_ne;  // fire, sampled on negedge

    always @(negedge clk)
        if (reset) fire_ne = 0; else fire_ne = fire;

    // Note:
    // - fire = [0, {{ntransitions-1}}] -> transition #fire is enabled
    // - fire = {{ntransitions}} -> all transitions are disabled

    fire_in_range : assume property ( `clk_rst fire <= {{ntransitions}} );

    fire_cycle_stable : assume property(`clk_rst fire == fire_ne);

    // model (derived from sg)

    integer state;

    always @(posedge clk or posedge reset) begin

        if (reset) begin

            {%- set initial_ind = state_inds[initial] %}

            state <= {{ initial_ind }}; // {{ initial }}

        end else begin
            {% for from, tr, to in transitions -%}
            {%- set signal = tr[:-1] -%}
            {%- set sign = tr[-1] -%}
            {%- set from_ind = state_inds[from] -%}
            {%- set to_ind = state_inds[to] -%}
            {%- set verilog_tr = ("~" + signal) if sign == "-" else signal %}
            if (state == {{ from_ind }} && {{ verilog_tr }} ) state <= {{ to_ind }};  // {{ to }}
            {%- endfor %}

        end

    end

    // Spec Compliance Properties:

    {%- for signal in inputs + outputs %}

    {%- set rise_tr = signal + "+" %}
    {%- set fall_tr = signal + "-" %}

    wire {{ signal }}_can_fall = 0
        {%- for prior, tr, _ in transitions if tr == fall_tr %}
        {%- set prior_ind = state_inds[prior] %}
        {{ "|| (state == %d)"|format(prior_ind) }}
        {%- endfor -%}
        ;

    wire {{ signal }}_can_rise = 0
        {%- for prior, tr, _ in transitions if tr == rise_tr %}
        {%- set prior_ind = state_inds[prior] %}
        {{ "|| (state == %d)"|format(prior_ind) }}
        {%- endfor -%}
        ;

    {%- endfor %}

    // Assumptions (spec compliance):
    {% for input in inputs %}
    compliance_{{input}}_rise: assume property ( `clk_rst $rose({{input}}) |-> {{input}}_can_rise );
    compliance_{{input}}_fall: assume property ( `clk_rst $fell({{input}}) |-> {{input}}_can_fall );
    {%- endfor %}

    // Assertions (spec compliance):
    {% for output in outputs %}
    compliance_{{output}}_rise: assert property ( `clk_rst $rose({{output}}) |-> {{output}}_can_rise );
    compliance_{{output}}_fall: assert property ( `clk_rst $fell({{output}}) |-> {{output}}_can_fall );
    {%- endfor %}

    // Enable signals:

    // Note: while internal transition enable status are indicated by (net ^
    // net_precap), inputs are generated by the environment and may therefore
    // may be enabled wile the expression (input ^ input_precap) is false.
    // Input enable status must therefore be derived from the spec, as
    // input_can_rise | input_can_fall.
    {% for input in inputs %}
    assign {{input}}_ena = {{input}}_can_rise | {{input}}_can_fall;
    {%- endfor -%}
    {%- for gate in stateful.values() %}
    {%- set output_net = get_output_net(gate) %}
    assign {{output_net}}_ena = {{output_net}}_precap ^ {{output_net}};
    {%- endfor %}

    // Output Persistency Properties:
    {% for gate in stateful.values() -%}
    {%- set output_net = get_output_net(gate) %}
    persistency_{{output_net}}: assert property ( `clk_rst {{output_net}}_ena |=> ({{output_net}}_ena || ~$stable({{output_net}})) );
    {%- endfor %}

    // Deadlock

    // Deadlock freeness: on each cycle, at least one internal transition is
    // enabled or an input can change.

    assign exist_enabled_transition =
        {%- for input in inputs %}
        | {{input}}_ena
        {%- endfor -%}
        {%- for gate in stateful.values() %}
        | {{ get_output_net(gate) }}_ena
        {%- endfor -%}
    ;

    // For arbiter circuit:
    //
    // always_grant: assert property ( `clk_rst
    //     $rose(r1) |-> ##[1:$] ($rose(g1) | $rose(g2) | $rose(g3) | exist_enabled_transition)
    // );

    deadlock_free: assert property ( `clk_rst
        not (##[1:$] ~exist_enabled_transition)
    );

    // Transition firing assumptions: a transitions can only be fired when
    // it's enabled (i.e. when a stateful gate can capture a new value = its
    // input and output are different).

    {% for input in inputs %}
    {%- set pre_net = input + "_precap" %}
    {%- set fire_ind = loop.index0 -%}
    firing_{{fire_ind}} : assume property ( `clk_rst (fire == {{fire_ind}}) |-> ({{input}} ^ {{pre_net}}) );
    {% endfor -%}

    {% for gate in stateful.values() %}
    {%- set output_net = get_output_net(gate) -%}
    {%- set pre_net = output_net + "_precap" %}
    {%- set fire_ind = loop.index0 + inputs|length -%}
    firing_{{fire_ind}} : assume property ( `clk_rst (fire == {{fire_ind}}) |-> ({{output_net}} ^ {{pre_net}}) );
    {% endfor %}
endmodule

module bind_info();

    bind circuit spec u1 (
          .reset(reset)
        , .clk(clk)
        , .fire(fire)

        {%- for input in inputs %}
        , .{{input}}({{ input }})
        , .{{input}}_precap({{ input }}_precap)
        {%- endfor %}

        {%- for gate in stateful.values() %}
        , .{{ get_output_net(gate) }}({{ get_output_net(gate) }})
        , .{{ get_output_net(gate) }}_precap({{ get_output_net(gate) }}_precap)
        {%- endfor -%}

    );

endmodule
