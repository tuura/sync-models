module Untitled (n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99);
    
    output n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;
    
    INV b0 (.I(n0), .ON(n1));
    BUF b1 (.I(n1), .O(n2));
    BUF b2 (.I(n2), .O(n3));
    BUF b3 (.I(n3), .O(n4));
    BUF b4 (.I(n4), .O(n5));
    BUF b5 (.I(n5), .O(n6));
    BUF b6 (.I(n6), .O(n7));
    BUF b7 (.I(n7), .O(n8));
    BUF b8 (.I(n8), .O(n9));
    BUF b9 (.I(n9), .O(n10));
    BUF b10 (.I(n10), .O(n11));
    BUF b11 (.I(n11), .O(n12));
    BUF b12 (.I(n12), .O(n13));
    BUF b13 (.I(n13), .O(n14));
    BUF b14 (.I(n14), .O(n15));
    BUF b15 (.I(n15), .O(n16));
    BUF b16 (.I(n16), .O(n17));
    BUF b17 (.I(n17), .O(n18));
    BUF b18 (.I(n18), .O(n19));
    BUF b19 (.I(n19), .O(n20));
    BUF b20 (.I(n20), .O(n21));
    BUF b21 (.I(n21), .O(n22));
    BUF b22 (.I(n22), .O(n23));
    BUF b23 (.I(n23), .O(n24));
    BUF b24 (.I(n24), .O(n25));
    BUF b25 (.I(n25), .O(n26));
    BUF b26 (.I(n26), .O(n27));
    BUF b27 (.I(n27), .O(n28));
    BUF b28 (.I(n28), .O(n29));
    BUF b29 (.I(n29), .O(n30));
    BUF b30 (.I(n30), .O(n31));
    BUF b31 (.I(n31), .O(n32));
    BUF b32 (.I(n32), .O(n33));
    BUF b33 (.I(n33), .O(n34));
    BUF b34 (.I(n34), .O(n35));
    BUF b35 (.I(n35), .O(n36));
    BUF b36 (.I(n36), .O(n37));
    BUF b37 (.I(n37), .O(n38));
    BUF b38 (.I(n38), .O(n39));
    BUF b39 (.I(n39), .O(n40));
    BUF b40 (.I(n40), .O(n41));
    BUF b41 (.I(n41), .O(n42));
    BUF b42 (.I(n42), .O(n43));
    BUF b43 (.I(n43), .O(n44));
    BUF b44 (.I(n44), .O(n45));
    BUF b45 (.I(n45), .O(n46));
    BUF b46 (.I(n46), .O(n47));
    BUF b47 (.I(n47), .O(n48));
    BUF b48 (.I(n48), .O(n49));
    BUF b49 (.I(n49), .O(n50));
    BUF b50 (.I(n50), .O(n51));
    BUF b51 (.I(n51), .O(n52));
    BUF b52 (.I(n52), .O(n53));
    BUF b53 (.I(n53), .O(n54));
    BUF b54 (.I(n54), .O(n55));
    BUF b55 (.I(n55), .O(n56));
    BUF b56 (.I(n56), .O(n57));
    BUF b57 (.I(n57), .O(n58));
    BUF b58 (.I(n58), .O(n59));
    BUF b59 (.I(n59), .O(n60));
    BUF b60 (.I(n60), .O(n61));
    BUF b61 (.I(n61), .O(n62));
    BUF b62 (.I(n62), .O(n63));
    BUF b63 (.I(n63), .O(n64));
    BUF b64 (.I(n64), .O(n65));
    BUF b65 (.I(n65), .O(n66));
    BUF b66 (.I(n66), .O(n67));
    BUF b67 (.I(n67), .O(n68));
    BUF b68 (.I(n68), .O(n69));
    BUF b69 (.I(n69), .O(n70));
    BUF b70 (.I(n70), .O(n71));
    BUF b71 (.I(n71), .O(n72));
    BUF b72 (.I(n72), .O(n73));
    BUF b73 (.I(n73), .O(n74));
    BUF b74 (.I(n74), .O(n75));
    BUF b75 (.I(n75), .O(n76));
    BUF b76 (.I(n76), .O(n77));
    BUF b77 (.I(n77), .O(n78));
    BUF b78 (.I(n78), .O(n79));
    BUF b79 (.I(n79), .O(n80));
    BUF b80 (.I(n80), .O(n81));
    BUF b81 (.I(n81), .O(n82));
    BUF b82 (.I(n82), .O(n83));
    BUF b83 (.I(n83), .O(n84));
    BUF b84 (.I(n84), .O(n85));
    BUF b85 (.I(n85), .O(n86));
    BUF b86 (.I(n86), .O(n87));
    BUF b87 (.I(n87), .O(n88));
    BUF b88 (.I(n88), .O(n89));
    BUF b89 (.I(n89), .O(n90));
    BUF b90 (.I(n90), .O(n91));
    BUF b91 (.I(n91), .O(n92));
    BUF b92 (.I(n92), .O(n93));
    BUF b93 (.I(n93), .O(n94));
    BUF b94 (.I(n94), .O(n95));
    BUF b95 (.I(n95), .O(n96));
    BUF b96 (.I(n96), .O(n97));
    BUF b97 (.I(n97), .O(n98));
    BUF b98 (.I(n98), .O(n99));
    BUF b99 (.I(n99), .O(n0));
    
    // signal values at the initial state:
    // !n0 !n1 !n2 !n3 !n4 !n5 !n6 !n7 !n8 !n9 !n10 !n11 !n12 !n13 !n14 !n15 !n16 !n17 !n18 !n19 !n20 !n21 !n22 !n23 !n24 !n25 !n26 !n27 !n28 !n29 !n30 !n31 !n32 !n33 !n34 !n35 !n36 !n37 !n38 !n39 !n40 !n41 !n42 !n43 !n44 !n45 !n46 !n47 !n48 !n49 !n50 !n51 !n52 !n53 !n54 !n55 !n56 !n57 !n58 !n59 !n60 !n61 !n62 !n63 !n64 !n65 !n66 !n67 !n68 !n69 !n70 !n71 !n72 !n73 !n74 !n75 !n76 !n77 !n78 !n79 !n80 !n81 !n82 !n83 !n84 !n85 !n86 !n87 !n88 !n89 !n90 !n91 !n92 !n93 !n94 !n95 !n96 !n97 !n98 !n99
    
endmodule
